`timescale 1ns/1ns

module DataPath_TB();

reg clk_tb;

DataPath uut(
    .clock(clk_tb));

initial begin
	$dumpfile("DataPath_TB.vcd");
    	$dumpvars(0, DataPath_TB);

	//Momento Ctrl + C & Ctrl + V

    	#100;
    	clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;

		clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
		clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	clk_tb = 1'b1;
    	#100;
        clk_tb = 1'b0;
    	#100;
    	
	
	$stop;
end   
endmodule


